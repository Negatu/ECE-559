framemem_inst : framemem PORT MAP (
		aclr	 => aclr_sig,
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
