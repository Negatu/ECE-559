library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;

entity FwdOutputCntrlr is
	port(clock,reset, dataRdEmpty, lengthRdEmpty : in std_logic; 
		 inFrameLengthValue: in std_logic_vector(20 downto 0);--11 bit length value + valid fram bit + 9 bit sequence number
		 lengthBuffer_RE,  dataBuffer_RE, fwdFrameValid: out std_logic;
		 fwdFrameLengthValue: out std_logic_vector(10 downto 0);
		 fwdSequenceNumbr : out std_logic_vector (8 downto 0));
end FwdOutputCntrlr;

architecture RegCountArch of FwdOutputCntrlr is
	
	component lengthValidReg IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (20 DOWNTO 0);
		enable		: IN STD_LOGIC ;
		q		    : OUT STD_LOGIC_VECTOR (20 DOWNTO 0)
	);
    END component;

	component outFrameLengthCounter IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		sclr		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (10 DOWNTO 0)
	);
   END component;
   
   component frameLengthValueComp IS
	PORT
	(
		dataa		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		AeB		    : OUT STD_LOGIC 
	);
    END component;
    	
	TYPE State_type IS ( NotEqual, Equal, RegWrite);
	SIGNAL y_current, y_next : State_type;
	signal counter_reset_sig, clear_length_reg, int_lengthBufferRE, equal_true, length_reg_we : std_logic; -- used to clear the counter after each frame
	signal int_FrameLengthValue : std_logic_vector(20 downto 0);
	signal counterValue : std_logic_vector (10 downto 0);
	
	begin
	
	lengthValidReg_inst : lengthValidReg PORT MAP (
		    aclr		=>  reset or clear_length_reg,
		    clock		=> clock,
			data     	=> inFrameLengthValue,
			enable		=> length_reg_we,
			q           => int_FrameLengthValue
	
		);
	outFrameLengthCounter_inst : outFrameLengthCounter PORT MAP (
		clock	=> clock,
		sclr	=> counter_reset_sig,
		q		=> counterValue
	
	);
	
	frameLengthValueComp_inst : frameLengthValueComp PORT MAP (
		dataa			=> int_FrameLengthValue (10 downto 0),
		datab			=> counterValue,
		AeB				=> equal_true
	);
	
	PROCESS(reset,clock)
	BEGIN
		IF Reset = '1' THEN y_current <= Equal;
		ELSIF clock'EVENT AND clock = '1' THEN
			y_current <= y_next;
		END IF;
	END PROCESS;
	
-- logic for determining next state
	PROCESS(dataRdEmpty, lengthRdEmpty, equal_true,y_current)
	BEGIN		
		CASE y_current IS
			WHEN NotEqual =>
				IF equal_true = '1' THEN y_next <= Equal;
				ELSE y_next <= NotEqual;
				END IF;
			WHEN Equal =>
				IF dataRdEmpty = '1' or lengthRdEmpty = '1' THEN y_next <= Equal;
				ELSE y_next <=  RegWrite;
				END IF;
			WHEN RegWrite =>
					y_next <= NotEqual;
		END CASE;
	END PROCESS;
	
-- output logic
	PROCESS(y_current, dataRdEmpty, lengthRdEmpty)
	BEGIN
		IF (y_current = Equal) THEN 
				dataBuffer_RE <= '0';
				counter_reset_sig <= '1';
				length_reg_we <= '0';
				IF dataRdEmpty = '1' or lengthRdEmpty = '1' THEN 
					int_lengthBufferRE <= '0';
					clear_length_reg <= '1';
				ELSE 
					int_lengthBufferRE <= '1';
					clear_length_reg <= '0';
				
				END IF;
				
				
		ELSIF (y_current = NotEqual) THEN
			dataBuffer_RE <= '1';
			int_lengthBufferRE <= '0';
			counter_reset_sig <= '0';
			clear_length_reg <= '0';
			length_reg_we <= '0';
		
		ELSE
			dataBuffer_RE <= '1';
			int_lengthBufferRE <= '0';
			counter_reset_sig <= '0';
			clear_length_reg <= '0';
			length_reg_we <= '1';
		
		END IF;
	END PROCESS;
	fwdFrameLengthValue <= int_FrameLengthValue(10 downto 0);
	fwdFrameValid		<= int_FrameLengthValue(11);
	fwdSequenceNumbr	<= int_frameLengthValue(20 downto 12);
	lengthBuffer_RE <= int_lengthBufferRE;
	
end RegCountArch;